module not_gate(
    ou,in
);
    input in;
    output ou;
    nand(ou,in,in);
endmodule 